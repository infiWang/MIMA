../def.sv