`include "def.sv"

module bubble (
    output reg [31:0] rdata
);

assign rdata = NOP;
    
endmodule