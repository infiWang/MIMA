enum bit [2:0] {
    f3OpInt_ADD = 3'b000,
    f3OpInt_AND = 3'b111,
    f3OpInt_OR = 3'b110,
    f3OpInt_XOR = 3'b100,
    f3OpInt_SL = 3'b001,
    f3OpInt_SR = 3'b101,
    f3OpInt_SLT = 3'b010,
    f3OpInt_SLTU = 3'b011
} f3OpInt;

enum bit [2:0] {
    f3Br_EQ = 3'b000,
    f3Br_NE = 3'b001,
    f3Br_LT = 3'b100,
    f3Br_GE = 3'b101,
    f3Br_LTU = 3'b110,
    f3Br_GEU = 3'b111
} f3Br;
