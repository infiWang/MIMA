../def.svh